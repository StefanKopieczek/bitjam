package color;
    typedef struct {
        logic [7:0] red;
        logic [7:0] green;
        logic [7:0] blue;        
    }  color_t;
endpackage